-- type generic for package
package p is
generic (
	type mytype
);
 
end package;