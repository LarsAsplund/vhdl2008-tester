-- this has to go wrong.
package t0 is
	big syntax error here
end package t0;
