-- ieee.fixed_generic_pkg
library ieee;
use ieee.fixed_generic_pkg.all;
package e9 is
end package e9;
