-- this can't go wrong.	
package t0 is
end package t0;
