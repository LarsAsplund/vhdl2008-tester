-- simple generic for package
package p is
generic (
	a:integer
);

end package;